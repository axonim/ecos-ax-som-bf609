# ====================================================================
#
#      i2c_lm3s.cdl
#
#      eCos Stellaris Cortex M3 I2C configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2011 Free Software Foundation, Inc.                        
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      ccoutand
# Contributors:
# Date:           2011-01-18
#
#####DESCRIPTIONEND####
# ====================================================================

cdl_package CYGPKG_DEVS_I2C_CORTEXM_LM3S {
    display       "I2C driver for Stellaris Cortex M3 microcontroller family"
    parent        CYGPKG_IO_I2C
    active_if     CYGPKG_IO_I2C
    active_if     CYGPKG_HAL_CORTEXM_LM3S
    include_dir   cyg/io
    description   "
        This package provides a generic I2C device driver for the on-chip
        I2C modules in Stellaris Cortex M3 microcontroller."

    compile       -library=libextras.a i2c_lm3s.c

    cdl_option CYGNUM_HAL_CORTEXM_LM3S_I2C_CLK_SPEED {
        display       "I2C channel clock"
        flavor        data
        default_value { 100000 }
        legal_values  { 100000 400000 }
        description   "
            Set the I2C clock speed. Slow mode (100KHz) or fast mode
            (400KHz)"
    }

    cdl_option CYGPKG_DEVS_I2C_CORTEXM_LM3S_TRACE {
        display       "I2C trace"
        flavor        bool
        default_value 0
        description   "
            Enable I2C transaction trace. Select to debug the driver."
    }

    cdl_component CYGPKG_DEVS_I2C_CORTEXM_LM3S_OPTIONS {
        display      "I2C driver build options"
        flavor        none
        active_if     { CYGINT_DEVS_I2C_CORTEXM_LM3S_BUS_DEVICES > 0 }
        description   "
            Package specific build options including control over
            compiler flags used only in building the Stellaris Cortex M3
            I2C bus driver."

        cdl_option CYGPKG_DEVS_I2C_CORTEXM_LM3S_CFLAGS_ADD {
            display       "Additional compiler flags"
            flavor        data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the Stellaris Cortex M3 I2C bus driver. These
                flags are used in addition to the set of global flags."
        }

        cdl_option CYGPKG_DEVS_I2C_CORTEXM_LM3S_CFLAGS_REMOVE {
            display       "Suppressed compiler flags"
            flavor        data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the Stellaris Cortex M3 I2C bus driver. These
                flags are removed from the set of global flags if
                present."
        }
    }
}

# EOF i2c_lm3s.cdl
