##=============================================================================
##
##      flash_m25pxx.cdl
##
##      M25Pxx SPI flash driver configuration options.
##
##=============================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2008, 2009 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
##=============================================================================
#######DESCRIPTIONBEGIN####
##
## Author(s):   Chris Holgate
## Date:        2008-12-22
## Purpose:     Configure M25Pxx SPI flash driver.
##
######DESCRIPTIONEND####
##
##=============================================================================

cdl_package CYGPKG_DEVS_FLASH_SPI_M25PXX {
    display	"M25PXX flash memory support"
    parent	CYGPKG_IO_FLASH
    active_if	CYGPKG_IO_FLASH CYGPKG_IO_SPI
    implements	CYGHWR_IO_FLASH_DEVICE
    implements  CYGHWR_IO_FLASH_INDIRECT_READS 
    include_dir	cyg/io
    compile	m25pxx.c

    description "
        Flash memory support for Numonyx M25Pxx SPI flash devices and 
        compatibles.  This driver implements the V2 flash driver API"

	cdl_option CYGNUM_DEVS_FLASH_SPI_M25PXX_READ_BLOCK_SIZE {
		display       "Maximum read block size"
		description   "
			In theory it is possible to read back the entire flash contents using
			a single SPI transaction.  However, some SPI bus drivers have a maximum 
			transaction size - for example transactions may be limited to the 
			length of a DMA bounce buffer.  Setting this option to a non-zero value 
			specifies the maximum SPI bus transfer size which will be used when 
			reading back data.  Read requests for areas larger than this block size 
			will automatically be split into a series of smaller SPI bus transactions.
		"
		flavor        data 
		default_value 0
	}
	

    cdl_option CYGPKG_DEVS_FLASH_SPI_M25PXX_TESTS {
        display "SPI Flash M25Pxx test"
        flavor  data
        calculated { "tests/m25pxx_test" }         
        description   "
            This option specifies the set of tests for the SPI m25pxx memory device drivers."
    }
}

# EOF flash_m25pxx.cdl