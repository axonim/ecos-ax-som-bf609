##==========================================================================
##
##      kinetis_fbram.cdl
##
##      Cortex-M Freescale Kinetis FBRAM configuration
##
##==========================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2010, 2011, 2012, 2013 Free Software Foundation, Inc.                  
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
##==========================================================================
#######DESCRIPTIONBEGIN####
##
## Author(s):    Ilija Kocho <ilijak@siva.com.mk>
## Date:         2013-04-28
##
######DESCRIPTIONEND####
##
##==========================================================================


#    cdl_component CYGPKG_HAL_CORTEXM_KINETIS_FBRAM {
#        display       "FlexBus RAM"
#        flavor bool
#        active_if     CYGINT_HAL_CORTEXM_KINETIS_DBRAM
#        default_value CYGINT_HAL_CORTEXM_KINETIS_FBRAM
#        description   "FlexBus RAM on Kinetis is mirrored at several address ranges.
#                Each mirror has its own caching options that may include:
#                non-cached, write-through and write-back.
#                By eCos configuration, FlexBus RAM is split in 3 partitions:
#                Cached, Non-cached and Code.
#                Cached partition is intended for general purpose main memory.
#                Non-cached partition is convenient for sharing
#                buffers with other bus masters such as Ethernet controller,
#                DMA, etc. Code partition is for executable code."
#

        cdl_option CYGHWR_HAL_KINETIS_FBR_SIZE {
            display       "FlexBus RAM size \[Bytes\]"
            flavor        data
            default_value CYGHWR_HAL_KINETIS_FB_CS0_SIZE ? CYGHWR_HAL_KINETIS_FB_CS0_SIZE * 1 : 0
        }

        cdl_option CYGHWR_HAL_KINETIS_FBR_SIZE_KIB {
            display       "FlexBus RAM size \[KiB\]"
            flavor        data
            calculated    { CYGHWR_HAL_KINETIS_FBR_SIZE / 1024 }
        }

        cdl_component CYGHWR_HAL_KINETIS_FBR_NON_CACHED_SIZE_KIB {
            display      "Non-cached FlexBus data RAM partition \[KiB\]"
            requires     { CYGHWR_HAL_KINETIS_FBR_NON_CACHED_SIZE_KIB <=
                           CYGHWR_HAL_KINETIS_FBR_SIZE_KIB }
            flavor       data

            implements   CYGINT_HAL_HAS_NONCACHED

            legal_values { 64 to (CYGHWR_HAL_KINETIS_FBR_SIZE_KIB - 64) }

            default_value { CYGHWR_HAL_KINETIS_FBR_SIZE_KIB / 4 }

            description "
                Non-cached FlexBus RAM partition, intended for sharing
                buffers with other bus masters such as Ethernet controller,
                DMA, etc."

            cdl_option CYGHWR_HAL_KINETIS_FBR_NON_CACHED_SIZE {
                display    "Non-cached FlexBus RAM size \[Bytes\]"
                flavor     data
                calculated { CYGHWR_HAL_KINETIS_FBR_NON_CACHED_SIZE_KIB
                             * 1024 * 0x1 }
            }

            cdl_option CYGHWR_HAL_KINETIS_FBR_NON_CACHED_BASE {
                display    "Non-cached FlexBus RAM base address"
                flavor     data

                calculated { CYGHWR_HAL_KINETIS_FBR_NON_CACHED_MIRROR +
                             CYGHWR_HAL_KINETIS_FBR_CACHED_SIZE +
                             CYGHWR_HAL_KINETIS_FBR_CODE_SIZE }
            }

            cdl_option CYGHWR_HAL_KINETIS_FBR_NON_CACHED_MIRROR {
                display       "Non-cached FlexBus RAM mirror base"
                flavor        data
                no_define
                legal_values     { 0x60000000 CYGINT_HAL_CORTEXM_KINETIS_150 ? 0x90000000 : 0x80000000 }
                default_value    { CYGINT_HAL_CORTEXM_KINETIS_150 ? 0x90000000 :
                                                                    0x60000000 }
            }

        }

        cdl_component CYGHWR_HAL_KINETIS_FBR_CODE_SIZE_KIB {
            display       "FlexBus RAM code partition \[KiB\]"
            requires      { CYGHWR_HAL_KINETIS_FBR_CODE_SIZE_KIB <=
                            CYGHWR_HAL_KINETIS_FBR_SIZE_KIB }
            flavor        data

            legal_values  { 64 to (CYGHWR_HAL_KINETIS_FBR_SIZE_KIB - 64) }

            default_value { CYGHWR_HAL_KINETIS_FBR_SIZE_KIB / 4 }

            description "
               FlexBus RAM code partition - for use as program memory.
               On systems with cache this partition is cached in PC cache
               and is always write-through"

            cdl_option CYGHWR_HAL_KINETIS_FBR_CODE_SIZE {
                display    "FlexBus RAM code partition size \[Bytes\]"
                flavor     data
                calculated { CYGHWR_HAL_KINETIS_FBR_CODE_SIZE_KIB
                             * 1024 * 0x1 }
            }

            cdl_option CYGHWR_HAL_KINETIS_FBR_CODE_BASE {
                display    "FlexBus RAM code partition base address"
                flavor     data

                legal_values     { 0x60000000
                                   CYGINT_HAL_CORTEXM_KINETIS_150 ? 0x18000000 :
                                                                    0x60000000 }
                default_value { CYGINT_HAL_CORTEXM_KINETIS_150 ? 0x18000000 :
                                                                 0x60000000 }
            }
        }

        cdl_component CYGHWR_HAL_KINETIS_FBR_CACHED_SIZE_KIB {
            display    "Cached FlexBus RAM data partition \[KiB\]"
            flavor     data
            requires   { CYGHWR_HAL_KINETIS_FBR_CACHED_SIZE_KIB >= 64 }
            calculated { CYGHWR_HAL_KINETIS_FBR_SIZE_KIB -
                         CYGHWR_HAL_KINETIS_FBR_NON_CACHED_SIZE_KIB -
                         CYGHWR_HAL_KINETIS_FBR_CODE_SIZE_KIB }

            description "
               Cached FlexBus RAM data partition - for general use as main data memory.
               On systems with cache this partition is cached in PS cache.
               Caching can be either copy-back or write-through and is determined
               by general cache mode setting."

            cdl_option CYGHWR_HAL_KINETIS_FBR_CACHED_SIZE {
                display    "Cached FlexBus RAM size \[Bytes\]"
                flavor      data
                calculated  { (CYGHWR_HAL_KINETIS_FBR_SIZE -
                              CYGHWR_HAL_KINETIS_FBR_NON_CACHED_SIZE -
                              CYGHWR_HAL_KINETIS_FBR_CODE_SIZE) * 0x1 }
                }

                cdl_option CYGHWR_HAL_KINETIS_FBR_CACHED_BASE {
                    display       "Cached FlexBus RAM base address"
                    flavor        data
                    calculated    { CYGHWR_HAL_KINETIS_FBR_CACHED_MIRROR +
                                    CYGHWR_HAL_KINETIS_FBR_CODE_SIZE }
                }

                cdl_option CYGHWR_HAL_KINETIS_FBR_CACHE_TYPE {
                    display     "FlexBus RAM cache type"
                    flavor       data
                    calculated  CYGSEM_HAL_DCACHE_STARTUP_MODE
                    description "FlexBus RAM cache type is determined by general
                        cache setting"
                }

                cdl_component CYGHWR_HAL_KINETIS_FBR_CACHED_MIRROR {
                    display         "Cached FlexBus RAM mirror base"
                    flavor data
                    no_define
                    legal_values     { 0x60000000 CYGINT_HAL_CORTEXM_KINETIS_150 ? 0x90000000 : 0x80000000 }
                    default_value    { 0x60000000 }
                    description      "Cached DDRAM base "
                }
        }

#    }

# EOF kinetis_fbram.cdl
