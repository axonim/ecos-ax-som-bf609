# ====================================================================
#
#      io_disk.cdl
#
#      eCos IO configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2003, 2009 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      savin
# Original data:  jskov, gthomas
# Contributors:
# Date:           2003-06-09
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_IO_DISK {
    display       "Disk device drivers"
    parent        CYGPKG_IO
    active_if     CYGPKG_IO
    requires      CYGPKG_ERROR
    include_dir   cyg/io
    description   "
        This option enables drivers for basic I/O services on
        disk devices."

    compile       -library=libextras.a disk.c
 
    define_proc {
        puts $::cdl_header "/***** proc output start *****/"
        puts $::cdl_header "#include <pkgconf/system.h>"
        puts $::cdl_header "#ifdef CYGDAT_IO_DISK_DEVICE_HEADER"
        puts $::cdl_header "# include CYGDAT_IO_DISK_DEVICE_HEADER"
        puts $::cdl_header "#endif "
        puts $::cdl_header "/****** proc output end ******/"
    }

    cdl_component CYGPKG_IO_DISK_DEVICES {
        display       "Hardware disk device drivers"
        flavor        bool
        default_value 1
        description   "
            This option enables the hardware disk drivers
            for the current platform."
    }

    cdl_component CYGDBG_IO_DISK_DEBUG {
        display       "Enable debugging output"
        flavor        bool
        default_value 0
        description   "
            This option enables debugging information from
            the disk driver package."
    }

    cdl_component CYGPKG_IO_DISK_OPTIONS {
        display "Disk device driver build options"
        flavor  none
        description   "
                Package specific build options including control over
                compiler flags used only in building this package,
                and details of which tests are built."


        cdl_option CYGPKG_IO_DISK_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the disk device drivers. These flags are used 
                in addition to the set of global flags."
        }

        cdl_option CYGPKG_IO_DISK_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the disk device drivers. These flags are removed from
                the set of global flags if present."
        }
    }
}

# ====================================================================
# EOF io_disk.cdl
