# ====================================================================
#
#      ser_cortexm_stm32.cdl
#
#      eCos serial ST STM32 configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2008, 2011 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      nickg
# Date:           2008-09-10
#
#####DESCRIPTIONEND####
#
# ====================================================================


cdl_package CYGPKG_IO_SERIAL_CORTEXM_STM32 {
    display       "ST STM32 serial device drivers"

    parent        CYGPKG_IO_SERIAL_DEVICES
    active_if     CYGPKG_IO_SERIAL
    active_if     CYGPKG_HAL_CORTEXM_STM32

    requires      CYGPKG_ERROR
    include_dir   cyg/io
    description   "
           This option enables the serial device drivers for the
           ST STM32."
    
    compile       -library=libextras.a   stm32_serial.c

    define_proc {
        puts $::cdl_system_header "/***** serial driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_DEVICE_HEADER <pkgconf/io_serial_cortexm_stm32.h>"
        puts $::cdl_system_header "/*****  serial driver proc output end  *****/"
    }

cdl_component CYGPKG_IO_SERIAL_CORTEXM_STM32_SERIAL0 {
    display       "ST STM32 serial port 0 driver"
    flavor        bool
    default_value CYGINT_HAL_STM32_UART0>0
    description   "
        This option includes the serial device driver for the ST STM32 
        port 0."

    cdl_option CYGDAT_IO_SERIAL_CORTEXM_STM32_SERIAL0_NAME {
        display       "Device name for ST STM32 serial port 0 driver"
        flavor        data
        default_value {"\"/dev/ser0\""}
        description   "
            This option specifies the name of the serial device for the 
            ST STM32 port 0."
    }

    cdl_option CYGNUM_IO_SERIAL_CORTEXM_STM32_SERIAL0_BAUD {
        display       "Baud rate for the ST STM32 serial port 0 driver"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 230400
        }
        default_value { CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD }
        description   "
            This option specifies the default baud rate (speed) for the 
            ST STM32 port 0."
    }

    cdl_option CYGNUM_IO_SERIAL_CORTEXM_STM32_SERIAL0_BUFSIZE {
        display       "Buffer size for the ST STM32 serial port 0 driver"
        flavor        data
        legal_values  0 to 8192
        default_value 128
        description   "
            This option specifies the size of the internal buffers used 
            for the ST STM32 port 0."
    }

    cdl_option CYGNUM_IO_SERIAL_CORTEXM_STM32_SERIAL0_INT_PRI {
        display       "Interrupt priority for STM32 serial port 0"
        flavor        data
        default_value 128
        legal_values  0 to 255
    }
}

cdl_component CYGPKG_IO_SERIAL_CORTEXM_STM32_SERIAL1 {
    display       "ST STM32 serial port 1 driver"
    flavor        bool
    default_value CYGINT_HAL_STM32_UART1>0
    description   "
        This option includes the serial device driver for the ST STM32 
        port 1."

    cdl_option CYGDAT_IO_SERIAL_CORTEXM_STM32_SERIAL1_NAME {
        display       "Device name for ST STM32 serial port 1 driver"
        flavor        data
        default_value {"\"/dev/ser1\""}
        description   "
            This option specifies the name of the serial device for the 
            ST STM32 port 1."
    }

    cdl_option CYGNUM_IO_SERIAL_CORTEXM_STM32_SERIAL1_BAUD {
        display       "Baud rate for the ST STM32 serial port 1 driver"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 230400
        }
        default_value CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD
        description   "
            This option specifies the default baud rate (speed) for the
            ST STM32 port 1."
    }

    cdl_option CYGNUM_IO_SERIAL_CORTEXM_STM32_SERIAL1_BUFSIZE {
        display       "Buffer size for the ST STM32 serial port 1 driver"
        flavor        data
        legal_values  0 to 8192
        default_value 128
        description   "
            This option specifies the size of the internal buffers used 
            for the ST STM32 port 1."
    }

    cdl_option CYGNUM_IO_SERIAL_CORTEXM_STM32_SERIAL1_INT_PRI {
        display       "Interrupt priority for STM32 serial port 1"
        flavor        data
        default_value 128
        legal_values  0 to 255
    }
}

cdl_component CYGPKG_IO_SERIAL_CORTEXM_STM32_SERIAL2 {
    display       "ST STM32 serial port 2 driver"
    flavor        bool
    default_value CYGINT_HAL_STM32_UART2>0
    description   "
        This option includes the serial device driver for the ST STM32 
        port 2."

    cdl_option CYGDAT_IO_SERIAL_CORTEXM_STM32_SERIAL2_NAME {
        display       "Device name for ST STM32 serial port 2 driver"
        flavor        data
        default_value {"\"/dev/ser2\""}
        description   "
            This option specifies the name of the serial device for the 
            ST STM32 port 2."
    }

    cdl_option CYGNUM_IO_SERIAL_CORTEXM_STM32_SERIAL2_BAUD {
        display       "Baud rate for the ST STM32 serial port 2 driver"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 230400
        }
        default_value CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD
        description   "
            This option specifies the default baud rate (speed) for the
            ST STM32 port 2."
    }

    cdl_option CYGNUM_IO_SERIAL_CORTEXM_STM32_SERIAL2_BUFSIZE {
        display       "Buffer size for the ST STM32 serial port 2 driver"
        flavor        data
        legal_values  0 to 8192
        default_value 128
        description   "
            This option specifies the size of the internal buffers used 
            for the ST STM32 port 2."
    }

    cdl_option CYGNUM_IO_SERIAL_CORTEXM_STM32_SERIAL2_INT_PRI {
        display       "Interrupt priority for STM32 serial port 2"
        flavor        data
        default_value 128
        legal_values  0 to 255
    }
}

cdl_component CYGPKG_IO_SERIAL_CORTEXM_STM32_SERIAL3 {
    display       "ST STM32 serial port 3 driver"
    flavor        bool
    default_value CYGINT_HAL_STM32_UART3>0
    description   "
        This option includes the serial device driver for the ST STM32 
        port 3."

    cdl_option CYGDAT_IO_SERIAL_CORTEXM_STM32_SERIAL3_NAME {
        display       "Device name for ST STM32 serial port 3 driver"
        flavor        data
        default_value {"\"/dev/ser3\""}
        description   "
            This option specifies the name of the serial device for the 
            ST STM32 port 3."
    }

    cdl_option CYGNUM_IO_SERIAL_CORTEXM_STM32_SERIAL3_BAUD {
        display       "Baud rate for the ST STM32 serial port 3 driver"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 230400
        }
        default_value CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD
        description   "
            This option specifies the default baud rate (speed) for the
            ST STM32 port 3."
    }

    cdl_option CYGNUM_IO_SERIAL_CORTEXM_STM32_SERIAL3_BUFSIZE {
        display       "Buffer size for the ST STM32 serial port 3 driver"
        flavor        data
        legal_values  0 to 8192
        default_value 128
        description   "
            This option specifies the size of the internal buffers used 
            for the ST STM32 port 3."
    }

    cdl_option CYGNUM_IO_SERIAL_CORTEXM_STM32_SERIAL3_INT_PRI {
        display       "Interrupt priority for STM32 serial port 3"
        flavor        data
        default_value 128
        legal_values  0 to 255
    }
}

cdl_component CYGPKG_IO_SERIAL_CORTEXM_STM32_SERIAL4 {
    display       "ST STM32 serial port 4 driver"
    flavor        bool
    default_value CYGINT_HAL_STM32_UART4>0
    description   "
        This option includes the serial device driver for the ST STM32 
        port 4."

    cdl_option CYGDAT_IO_SERIAL_CORTEXM_STM32_SERIAL4_NAME {
        display       "Device name for ST STM32 serial port 4 driver"
        flavor        data
        default_value {"\"/dev/ser4\""}
        description   "
            This option specifies the name of the serial device for the 
            ST STM32 port 4."
    }

    cdl_option CYGNUM_IO_SERIAL_CORTEXM_STM32_SERIAL4_BAUD {
        display       "Baud rate for the ST STM32 serial port 4 driver"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 230400
        }
        default_value CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD
        description   "
            This option specifies the default baud rate (speed) for the
            ST STM32 port 4."
    }

    cdl_option CYGNUM_IO_SERIAL_CORTEXM_STM32_SERIAL4_BUFSIZE {
        display       "Buffer size for the ST STM32 serial port 4 driver"
        flavor        data
        legal_values  0 to 8192
        default_value 128
        description   "
            This option specifies the size of the internal buffers used 
            for the ST STM32 port 4."
    }

    cdl_option CYGNUM_IO_SERIAL_CORTEXM_STM32_SERIAL4_INT_PRI {
        display       "Interrupt priority for STM32 serial port 4"
        flavor        data
        default_value 128
        legal_values  0 to 255
    }
}

cdl_component CYGPKG_IO_SERIAL_CORTEXM_STM32_SERIAL5 {
    display       "ST STM32 serial port 5 driver"
    flavor        bool
    default_value CYGINT_HAL_STM32_UART5>0
    description   "
        This option includes the serial device driver for the ST STM32 
        port 5."

    cdl_option CYGDAT_IO_SERIAL_CORTEXM_STM32_SERIAL5_NAME {
        display       "Device name for ST STM32 serial port 5 driver"
        flavor        data
        default_value {"\"/dev/ser5\""}
        description   "
            This option specifies the name of the serial device for the 
            ST STM32 port 5."
    }

    cdl_option CYGNUM_IO_SERIAL_CORTEXM_STM32_SERIAL5_BAUD {
        display       "Baud rate for the ST STM32 serial port 5 driver"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 230400
        }
        default_value CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD
        description   "
            This option specifies the default baud rate (speed) for the
            ST STM32 port 5."
    }

    cdl_option CYGNUM_IO_SERIAL_CORTEXM_STM32_SERIAL5_BUFSIZE {
        display       "Buffer size for the ST STM32 serial port 5 driver"
        flavor        data
        legal_values  0 to 8192
        default_value 128
        description   "
            This option specifies the size of the internal buffers used 
            for the ST STM32 port 5."
    }

    cdl_option CYGNUM_IO_SERIAL_CORTEXM_STM32_SERIAL5_INT_PRI {
        display       "Interrupt priority for STM32 serial port 5"
        flavor        data
        default_value 128
        legal_values  0 to 255
    }
}


    cdl_component CYGPKG_IO_SERIAL_CORTEXM_STM32_OPTIONS {
        display "Serial device driver build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_IO_SERIAL_CORTEXM_STM32_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_IO_SERIAL_CORTEXM_STM32_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are removed from
                the set of global flags if present."
        }
    }

    cdl_component CYGPKG_IO_SERIAL_CORTEXM_STM32_TESTING {
        display    "Testing parameters"
        flavor     none

        implements CYGINT_IO_SERIAL_TEST_SKIP_115200
        implements CYGINT_IO_SERIAL_TEST_SKIP_57600
        implements CYGINT_IO_SERIAL_TEST_SKIP_38400

        cdl_option CYGPRI_SER_TEST_SER_DEV {
            display       "Serial device used for testing"
            flavor        data
            default_value { CYGPKG_IO_SERIAL_CORTEXM_STM32_SERIAL0 ? CYGDAT_IO_SERIAL_CORTEXM_STM32_SERIAL0_NAME : \
                            CYGPKG_IO_SERIAL_CORTEXM_STM32_SERIAL1 ? CYGDAT_IO_SERIAL_CORTEXM_STM32_SERIAL1_NAME : \
                            CYGPKG_IO_SERIAL_CORTEXM_STM32_SERIAL2 ? CYGDAT_IO_SERIAL_CORTEXM_STM32_SERIAL2_NAME : \
                            CYGPKG_IO_SERIAL_CORTEXM_STM32_SERIAL3 ? CYGDAT_IO_SERIAL_CORTEXM_STM32_SERIAL3_NAME : \
                            CYGPKG_IO_SERIAL_CORTEXM_STM32_SERIAL4 ? CYGDAT_IO_SERIAL_CORTEXM_STM32_SERIAL4_NAME : \
                            CYGDAT_IO_SERIAL_CORTEXM_STM32_SERIAL5_NAME }
        }

        cdl_option CYGPRI_SER_TEST_TTY_DEV {
            display       "TTY-mode serial device used for testing"
            flavor        data
            default_value { CYGPKG_IO_SERIAL_CORTEXM_STM32_SERIAL0 ? "\"/dev/tty0\"" : \
                            CYGPKG_IO_SERIAL_CORTEXM_STM32_SERIAL1 ? "\"/dev/tty1\"" : \
                            CYGPKG_IO_SERIAL_CORTEXM_STM32_SERIAL2 ? "\"/dev/tty2\"" : \
                            CYGPKG_IO_SERIAL_CORTEXM_STM32_SERIAL3 ? "\"/dev/tty3\"" : \
                            CYGPKG_IO_SERIAL_CORTEXM_STM32_SERIAL4 ? "\"/dev/tty4\"" : \
                            "\"/dev/tty5\"" }
        }

        define_proc {
            puts $::cdl_header "#define CYGPRI_SER_TEST_CRASH_ID \"stm32\""
        }
    }
}

# EOF ser_cortexm_stm32.cdl
