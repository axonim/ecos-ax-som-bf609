# ====================================================================
#
#      devs_flash_atmel_dataflash.cdl
#
#      Atmel DataFlash parts support
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Savin Zlobec <savin@elatec.si> 
# Date:           2004-08-27
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_FLASH_ATMEL_DATAFLASH {
    display       "Atmel DataFlash parts support"
    description   "Support for Atmel DataFlash"
    parent        CYGPKG_IO_FLASH
    active_if	  CYGPKG_IO_SPI
    requires      CYGPKG_ERROR    
    hardware
    compile       devs_flash_atmel_dataflash.c 
    include_dir   cyg/io

    cdl_interface CYGPKG_DEVS_FLASH_ATMEL_DATAFLASH_FLASH_DEV {
        display         "Support for DataFlash IO Flash interface"
        flavor          bool
        active_if       CYGPKG_IO_FLASH
        implements      CYGHWR_IO_FLASH_DEVICE
	implements	CYGHWR_IO_FLASH_INDIRECT_READS
        compile         devs_flash_atmel_dataflash_flash_dev_funs.c     
        description     "This option will be enabled by platforms which
            need to support access to DataFlash through IO Flash API."
    }
}

# EOF devs_flash_atmel_dataflash.cdl 
