# ====================================================================
#
#      ser_MCF5272_uart.cdl
#
#      eCos serial driver for MCF5272 UART
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2006 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================

cdl_package CYGPKG_IO_SERIAL_COLDFIRE_MCF5272 {
    display       "Serial driver for MCF5272 UART"

    parent        CYGPKG_IO_SERIAL_DEVICES
    active_if     CYGPKG_IO_SERIAL
    requires      CYGPKG_ERROR
    include_dir   cyg/io
    description   "
           This option enables the serial device drivers for the
           ColdFire MCF5272."

    compile       -library=libextras.a mcf5272_serial.c

    cdl_component CYGPKG_IO_SERIAL_COLDFIRE_MCF5272_CHANNEL0 {
        display       "MCF5272 UART serial port 0 driver"
        flavor        bool
        default_value 1

        implements    CYGINT_IO_SERIAL_FLOW_CONTROL_HW
        implements    CYGINT_IO_SERIAL_LINE_STATUS_HW

        description   "This option includes the serial device driver
            for the MCF5272 UART port 0."

        cdl_option CYGDAT_IO_SERIAL_COLDFIRE_MCF5272_CHANNEL0_NAME {
            display       "Device name for the MCF5272 UART serial port 0"
            flavor        data
            default_value {"\"/dev/ser0\""}
            description   "
                This option specifies the name of serial device for the
                MCF5272 UART port 0."
         }

        cdl_option CYGNUM_IO_SERIAL_COLDFIRE_MCF5272_CHANNEL0_BAUD {
            display       "Baud rate for the MCF5272 UART serial port 0"
            flavor        data
            legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                          4800 7200 9600 14400 19200 38400 57600 115200 230400
            }
            default_value 19200
            description   "
                This option specifies the default baud rate (speed) for the
                MCF5272 UART port 0."
        }

        cdl_option CYGOPT_IO_SERIAL_COLDFIRE_MCF5272_CHANNEL0_AUTOBAUD {
            display       "Enable automatic baud rate detection for the MCF5272 UART serial port 0."
            flavor        bool
            default_value 0
            active_if     CYGNUM_IO_SERIAL_COLDFIRE_MCF5272_CHANNEL0_BUFSIZE > 0
            description   "
                This option enables automatic baud rate detection for
                MCF5272 UART port 0. Sending a BREAK character on the
                line will start the detection. The first character following
                the BREAK should occupy an odd position in the character table
                (like \'a\'). This option requires interrupts to be enabled
                for the port."
        }

        cdl_option CYGNUM_IO_SERIAL_COLDFIRE_MCF5272_CHANNEL0_BUFSIZE {
            display       "Buffer size for the MCF5272 UART serial port 0"
            flavor        data
            legal_values  0 to 8192
            default_value 128
            description   "
                This option specifies the size of the internal buffers used
                for the MCF5272 UART port 0. If the size specified is 0, the
                driver will not use interrupts."
        }

        cdl_option CYGNUM_IO_SERIAL_COLDFIRE_MCF5272_CHANNEL0_PRIORITY {
            display       "Interrupt priority level for MCF5272 UART serial port 0"
            flavor        data
            legal_values  1 to 6
            default_value 2
            active_if     CYGNUM_IO_SERIAL_COLDFIRE_MCF5272_CHANNEL0_BUFSIZE > 0
            description   "
                This option specifies the priority associated to interrupts
                coming from the MCF5272 UART port 0."
        }
    }

    cdl_component CYGPKG_IO_SERIAL_COLDFIRE_MCF5272_CHANNEL1 {
        display       "MCF5272 UART serial port 1 driver"
        flavor        bool
        default_value 0

        implements    CYGINT_IO_SERIAL_FLOW_CONTROL_HW
        implements    CYGINT_IO_SERIAL_LINE_STATUS_HW

        description   "This option includes the serial device driver for the
            MCF5272 UART port 1."

        cdl_option CYGDAT_IO_SERIAL_COLDFIRE_MCF5272_CHANNEL1_NAME {
            display       "Device name for the MCF5272 UART serial port 1"
            flavor        data
            default_value {"\"/dev/ser1\""}
            description   "
                This option specifies the name of serial device for the
                MCF5272 UART port 1."
         }

        cdl_option CYGNUM_IO_SERIAL_COLDFIRE_MCF5272_CHANNEL1_BAUD {
            display       "Baud rate for the MCF5272 UART serial port 1"
            flavor        data
            legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                          4800 7200 9600 14400 19200 38400 57600 115200 230400
            }
            default_value 19200
            description   "
                This option specifies the default baud rate (speed) for the
                MCF5272 UART port 1."
        }

        cdl_option CYGOPT_IO_SERIAL_COLDFIRE_MCF5272_CHANNEL1_AUTOBAUD {
            display       "Enable automatic baud rate detection for the MCF5272 UART serial port 1."
            flavor        bool
            default_value 0
            active_if     CYGNUM_IO_SERIAL_COLDFIRE_MCF5272_CHANNEL1_BUFSIZE > 0
            description   "
                This option enables automatic baud rate detection for
                MCF5272 UART port 1. Sending a BREAK character on the
                line will start the detection. The first character following
                the BREAK should occupy an odd position in the character table
                (like \'a\'). This option requires interrupts to be enabled
                for the port."
        }

        cdl_option CYGNUM_IO_SERIAL_COLDFIRE_MCF5272_CHANNEL1_BUFSIZE {
            display       "Buffer size for the MCF5272 UART serial port 1"
            flavor        data
            legal_values  0 to 8192
            default_value 128
            description   "
                This option specifies the size of the internal buffers used
                for the MCF5272 UART port 1. If the size specified is 0, the
                driver will not use interrupts."
        }

        cdl_option CYGNUM_IO_SERIAL_COLDFIRE_MCF5272_CHANNEL1_PRIORITY {
            display       "Interrupt priority level for MCF5272 UART serial port 1"
            flavor        data
            legal_values  1 to 6
            default_value 2
            active_if     CYGNUM_IO_SERIAL_COLDFIRE_MCF5272_CHANNEL1_BUFSIZE > 0
            description   "
                This option specifies the priority associated to interrupts
                coming from the MCF5272 UART port 1."
        }
    }
}

