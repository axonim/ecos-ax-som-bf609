# ====================================================================
#
#      i2c_a2fxxx.cdl
#
#      eCos Smartfusion Cortex-M3 I2C configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2011 Free Software Foundation, Inc.                        
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      ccoutand
# Contributors:
# Date:           2011-01-18
#
#####DESCRIPTIONEND####
# ====================================================================

cdl_package CYGPKG_DEVS_I2C_CORTEXM_A2FXXX  {
    display       "Actel Smartfusion I2C driver"
    parent        CYGPKG_IO_I2C
    active_if     CYGPKG_IO_I2C
    active_if     CYGPKG_HAL_CORTEXM_A2FXXX
    include_dir   cyg/io
    description   "
        This package provides a generic I2C device driver for the on-chip
        I2C modules in Smartfusion Cortex-M3 microcontroller."

    compile       -library=libextras.a i2c_a2fxxx.c

    cdl_option CYGNUM_HAL_CORTEXM_A2FXXX_I2C_CLK_DIV {
        display       "I2C channel clock divider"
        flavor        data
        default_value { 256 }
        legal_values  { 8 60 120 160 192 960 224 256 960}
        description   "
            Set the I2C clock divider."
    }

    cdl_option CYGDBG_DEVS_I2C_CORTEXM_A2FXXX_TRACE {
        display       "Display status messages during I2C operations"
        flavor        bool
        default_value 0
        description   "
           Selecting this option will cause the I2C driver to print status
           messages as various I2C operations are undertaken."
    }

    cdl_component CYGPKG_DEVS_I2C_CORTEXM_A2FXXX_OPTIONS {
        display      "I2C driver build options"
        flavor        none
        active_if     { CYGINT_DEVS_I2C_CORTEXM_A2FXXX_BUS_DEVICES > 0 }
        description   "
            Package specific build options including control over
            compiler flags used only in building the Smartfusion Cortex-M3
            I2C bus driver."

        cdl_option CYGPKG_DEVS_I2C_CORTEXM_A2FXXX_CFLAGS_ADD {
            display       "Additional compiler flags"
            flavor        data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the Smartfusion Cortex-M3 I2C bus driver. These
                flags are used in addition to the set of global flags."
        }

        cdl_option CYGPKG_DEVS_I2C_CORTEXM_A2FXXX_CFLAGS_REMOVE {
            display       "Suppressed compiler flags"
            flavor        data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the Smartfusion Cortex-M3 I2C bus driver. These
                flags are removed from the set of global flags if
                present."
        }
    }
}

# EOF i2c_a2fxxx.cdl
