# ====================================================================
#
#      ser_loop.cdl
#
#      eCos serial LOOP configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2009 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  gthomas
# Contributors:
# Date:           1999-07-07
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_IO_SERIAL_LOOP {
    display       "Loop serial device drivers"

    parent        CYGPKG_IO_SERIAL_DEVICES
    active_if     CYGPKG_IO_SERIAL
    requires      CYGPKG_ERROR
    include_dir   cyg/io
    include_files ; # none _exported_ whatsoever

    description   "
       This package contains the loop serial device driver."

    compile       -library=libextras.a loop_serial.c

    # FIXME: Bad name
    cdl_option CYGPKG_IO_SERIAL_LOOP_POLLED_MODE {
        display       "LOOP polled mode serial drivers"
        flavor        bool
        default_value 0
        description   "
            If asserted, this option specifies that the serial loop device
            drivers for the should be polled-mode instead of
            interrupt driven."
    }
    
    cdl_component CYGPKG_IO_SERIAL_LOOP_SERIAL0 {
        display       "LOOP serial port 0 driver"
        flavor        bool
        default_value 0
        description   "
            This option includes the serial loop device driver for port 0." 
    
        cdl_option CYGDAT_IO_SERIAL_LOOP_SERIAL0_NAME {
            display       "Device name for LOOP serial port 0"
            flavor        data
            default_value {"\"/dev/ser0\""}
            description   "
                This option specifies the first loop device name."
        }
    
        cdl_option CYGNUM_IO_SERIAL_LOOP_SERIAL0_BAUD {
            display       "Baud rate for the LOOP serial port 0 driver"
            flavor        data
            legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800
                            2400 3600 4800 7200 9600 14400 19200 38400
                            57600 115200 230400
            }
            default_value 38400
            description   "
                This option specifies the default baud rate (speed) for the
                LOOP port 0."
        }
    
        cdl_option CYGNUM_IO_SERIAL_LOOP_SERIAL0_BUFSIZE {
            display       "Buffer size for the LOOP serial port 0 driver"
            flavor        data
            legal_values  0 to 8192
            default_value 128
            description   "
                This option specifies the size of the internal buffers used
                for the LOOP port 0."
        }
    }
    
    cdl_component CYGPKG_IO_SERIAL_LOOP_SERIAL1 {
        display       "LOOP serial port 1 driver"
        flavor        bool
        default_value 0
        description   "
            This option includes the serial device driver for port 1 on
            the LOOP."
    
        cdl_option CYGDAT_IO_SERIAL_LOOP_SERIAL1_NAME {
            display       "Device name for LOOP serial port 1"
            flavor        data
            default_value {"\"/dev/ser1\""}
            description   "
                This option specifies the device name port 1 on the LOOP."
        }
    
        cdl_option CYGNUM_IO_SERIAL_LOOP_SERIAL1_BAUD {
            display       "Baud rate for the LOOP serial port 1 driver"
            flavor        data
            legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800
                            2400 3600 4800 7200 9600 14400 19200 38400
                            57600 115200 230400
            }
            default_value 38400
            description   "
                This option specifies the default baud rate (speed) for the
                LOOP port 1."
        }
    
        cdl_option CYGNUM_IO_SERIAL_LOOP_SERIAL1_BUFSIZE {
            display       "Buffer size for the LOOP serial port 1 driver"
            flavor        data
            legal_values  0 to 8192
            default_value 128
            description   "
                This option specifies the size of the internal buffers used
                for the LOOP port 1."
        }
    }

    cdl_component CYGPKG_IO_SERIAL_LOOP_OPTIONS {
        display "Serial device driver build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_IO_SERIAL_LOOP_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags
                are used in addition to the set of global flags."
        }

        cdl_option CYGPKG_IO_SERIAL_LOOP_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are
                removed from the set of global flags if present."
        }
    }
}

# EOF ser_loop.cdl
