## ====================================================================
##
##      flash_stm32.cdl
##
##      FLASH memory - Hardware support for STM32 on-chip flash
##
## ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2008, 2011 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
## ====================================================================
######DESCRIPTIONBEGIN####
##
## Author(s):      nickg
## Date:           2008-09-22
##
#####DESCRIPTIONEND####
##
## ====================================================================

cdl_package CYGPKG_DEVS_FLASH_STM32 {
    display       "STM32 FLASH memory support"
    parent        CYGPKG_IO_FLASH
    active_if	  CYGPKG_IO_FLASH
    implements    CYGHWR_IO_FLASH_DEVICE

    include_dir   cyg/io

    compile	  stm32_flash.c

    description "
        Flash memory support for on-chip flash on STM32 devices and compatibles.
        This driver implements the V2 flash driver API."

    cdl_option CYGNUM_DEVS_FLASH_STM32_V2_PROGRAM_BURST_SIZE {
	display		"Number of words to write per burst"
	flavor		data
	default_value	256
	legal_values	4 to 4096
	description "
            On typical hardware programming the flash requires disabling
            interrupts for an extended period of time.
            Some or all of the flash hardware will be unusable while each word
            is programmed, and disabling interrupts is the only reliable
            way of ensuring that no interrupt handler or other thread will
            try to access the flash in the middle of an operation. This
            can have a major impact on the real-time responsiveness of
            typical applications. To ameliorate this the driver will
            perform writes in small bursts, briefly re-enabling the cache
            and interrupts between each burst. The number of write operations
            per burst is determined by this option: reducing the number of
            writes per burst will improve real-time response, but will add
            overhead so the actual flash program operation will take
            longer; conversely more writes per burst will worsen response
            times but reduce overhead."
    }
    
    cdl_option CYGNUM_DEVS_FLASH_STM32_PARALLELISM {
        display         "Program/erase parallelism"
        flavor          data
        legal_values    { 8 16 32 64 }
        active_if       { ((CYGHWR_HAL_CORTEXM_STM32_FAMILY == "F2") || (CYGHWR_HAL_CORTEXM_STM32_FAMILY == "F4")) }
        default_value   32
        description     "
            The Flash interface of the STM32 F2 and F4 families can program or erase
            multiple bits in one step. The maximum possible parallelism depends
            on the supply voltage. The default value of this option (32)
            corresponds to supply voltage of 2.7 - 3.6V, but another value
            may be chosen if a different voltage is used."
    }
    
    cdl_component CYGPKG_DEVS_FLASH_STM32_OPTIONS {
        display "STM32 driver build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building the STM32
            flash driver, and details of which tests are built."

        cdl_option CYGPKG_DEVS_FLASH_STM32_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the STM32 flash driver. These flags
                are used in addition to the set of global flags."
        }

        cdl_option CYGPKG_DEVS_FLASH_STM32_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the STM32 flash driver. These flags
                are removed from the set of global flags if present."
        }
    }
}

# End of flash_stm32.cdl
