# ====================================================================
#
#      objloader.cdl
#
#      Object loader configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2005, 2008, 2009 Free Software Foundation, Inc.                        
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Anthony Tonizzo (atonizzo@gmail.com)
# Contributors:   Andrew Lunn
# Date:           2005-05-13
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_OBJLOADER {
    display       "Object file loader"
    description   "This package provides support for loading and relocating 
                   object files within eCos."
    include_dir   cyg/objloader
    include_files elf.h objelf.h loader_fs.h relocate_ppc.h relocate_i386.h
    include_files relocate_arm.h loader_memory.h
    compile       objloader.c objelf.c
    requires      CYGPKG_MEMALLOC
# ====================================================================

    cdl_component CYGPKG_SERVICES_OBJLOADER_ARCHITECTURE {
        display "Architecture dependent settings"
        flavor  none
        no_define
        requires CYGINT_SERVICES_OBJLOADER_RELOCATOR == 1

        description   "Each of the options here enables the correct
                       relocation support for the architectures supported."

        cdl_interface CYGINT_SERVICES_OBJLOADER_RELOCATOR {
            display "Suitable function to perform a symbol relocation"
            description "
                For each architecture we need a function which relocate
                a symbol. If we don't have a relocator the loader
                cannot work."
        }

        cdl_option CYGBLD_OBJLOADER_ARCHITECTURE_POWERPC {
           display       "Support loading on PowerPC processors"
           calculated    CYGPKG_HAL_POWERPC
           implements    CYGINT_SERVICES_OBJLOADER_RELOCATOR
           define_proc {
               puts $::cdl_header "#include <cyg/objloader/relocate_ppc.h>"
           }
           compile relocate_ppc.c
        }

        cdl_option CYGBLD_OBJLOADER_ARCHITECTURE_I386 {
           display       "Support loading on I386 processors"
           calculated    CYGPKG_HAL_I386 || CYGPKG_HAL_SYNTH_I386
           implements    CYGINT_SERVICES_OBJLOADER_RELOCATOR
           define_proc {
               puts $::cdl_header "#include <cyg/objloader/relocate_i386.h>"
           }
           compile relocate_i386.c
        }

        cdl_option CYGBLD_OBJLOADER_ARCHITECTURE_ARM {
            display       "Support loading on ARM processors"
            calculated    CYGPKG_HAL_ARM
            implements    CYGINT_SERVICES_OBJLOADER_RELOCATOR
            define_proc {
               puts $::cdl_header "#include <cyg/objloader/relocate_arm.h>"
            }
            compile relocate_arm.c
        }
        
    }
 
    cdl_component CYGOPT_SERVICES_OBJLOADER_LOADERS {
        display "Loaders to compile"
        flavor  none
        no_define
        description   "Options to select which types of loaders (e.g. from file
                       system, memory, http etc. to compile."

      cdl_option CYGOPT_SERVICES_OBJLOADER_LOADERS_FS {
          display       "Load module from file system"
          flavor        bool
          default_value 1
          requires      CYGPKG_IO_FILEIO
          description   "This option will compile the code required to load an
                         object library from a generic file system." 
          compile       loader_fs.c
      }

      cdl_option CYGOPT_SERVICES_OBJLOADER_LOADERS_MEMORY {
          display       "Load module from memory"
          flavor        bool
          default_value 1
          description   "This option will compile the module required to load an
                         object library from a ROM memory." 
          compile       loader_memory.c
      }
    }  

    cdl_option CYGPKG_SERVICES_OBJLOADER_DEBUG_LEVEL {
        display          "Verbosity of debug output"
        flavor           data
        legal_values     0 1 2
        default_value    0
        description      "This option allows controls over the verbosity of
                         the debug output. 1 is moderate, 2 is very
                         verbose, including the symbol name of each relocation
                         performed. Any value other than 0 will prevent the
                         unloading of unused library data, thus increasing the
                         heap memory requirements of the package."
    }
   
    cdl_component CYGPKG_SERVICES_OBJLOADER_OPTIONS {
        display "Object loader build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_SERVICES_OBJLOADER_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the serial device drivers. These flags are
                used in addition to the set of global flags."
        }

        cdl_option CYGPKG_SERVICES_OBJLOADER_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the serial device drivers. These flags are
                removed from the set of global flags if present."
        }
    }

    cdl_component CYGTST_SERVICES_OBJLOADER_BUILD_TESTS {
        display       "Build test library"
        default_value 0
        active_if     CYGPKG_FS_ROM
        active_if     CYGINT_SERVICES_OBJLOADER_RELOCATOR
        requires      CYGBLD_FS_ROMFS_MK_ROMFS
        no_define
        description   "
            This option enables the building of a library and an
            application for testing the loader." 
        
        make -priority 320 {
            testobj/hello.o : <PACKAGE>/tests/library/hello.c
            @mkdir -p "$(dir $@)"
            $(CC) -c $(INCLUDE_PATH) -I$(dir $<) $(ACTUAL_CFLAGS) -o $@ $<
        }

        make -priority 322 {
            <PREFIX>/include/cyg/objloader/testromfs_be.h : testobj/hello.o
            $(PREFIX)/bin/mk_romfs -b $(dir $<) testromfs_be.bin
            @mkdir -p "$(dir $@)"
            @tclsh $(PREFIX)/bin/file2c.tcl testromfs_be.bin $@
        }
        
        make -priority 322 {
            <PREFIX>/include/cyg/objloader/testromfs_le.h : testobj/hello.o
            $(PREFIX)/bin/mk_romfs $(dir $<) testromfs_le.bin
            @mkdir -p "$(dir $@)"
            @tclsh $(PREFIX)/bin/file2c.tcl testromfs_le.bin $@
        }
    
        cdl_option CYGPKG_OBJLOADER_TESTS {
            display     "Objloader tests"
            flavor      data
            no_define
            calculated  { "tests/test_mods" }
            description "
                This option specifies the set of tests for the object
                loader package"
       }
    }
}

# ====================================================================
# EOF objloader.cdl
