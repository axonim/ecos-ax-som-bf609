# ====================================================================
#
#      hal_arm_at91.cdl
#
#      Atmel AT91 HAL package configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2003, 2010 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Contributors:   gthomas, tkoeller, tdrury, nickg, jld
# Date:           2001-07-12
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_ARM_AT91 {
    display       "Atmel AT91 variant HAL"
    parent        CYGPKG_HAL_ARM
    define_header hal_arm_at91.h
    include_dir   cyg/hal
    hardware
    description   "
        The AT91 HAL package provides the support needed to run
        eCos on Atmel AT91 based targets."

    compile       at91_misc.c

    implements    CYGINT_HAL_DEBUG_GDB_STUBS
    implements    CYGINT_HAL_DEBUG_GDB_STUBS_BREAK
    implements    CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT
    implements    CYGINT_HAL_VIRTUAL_VECTOR_COMM_BAUD_SUPPORT
    implements    CYGINT_HAL_ARM_ARCH_ARM7
    implements    CYGINT_HAL_ARM_THUMB_ARCH

    # Let the architectural HAL see this variant's files
    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_ARM_VAR_IO_H"
        puts $::cdl_system_header "#define CYGBLD_HAL_ARM_VAR_ARCH_H"
    }

    cdl_option CYGHWR_HAL_ARM_AT91 {
        display        "AT91 variant used"
        flavor         data
        default_value  {"R40807"}
        legal_values   {"R40807" "R40008" "M42800A" "M55800A" "JTST" 
                        "AT91SAM7S" }
        description    "The AT91 microcontroller family has several variants,
                        the main differences being the amount of on-chip SRAM,
                        peripherals and their layout. This option allows the
                        platform HALs to select the specific microcontroller
                        being used."
    }

    cdl_option CYGHWR_HAL_ARM_AT91_FIQ {
        display       "handle FIQ as an IRQ"
        flavor        bool
        default_value 0
        description   "
            Enable this option if you need to handle FIQ interrupts in the
            normal way, i.e. a FIQ interrupt will be treated as a normal IRQ 
            using the highest priority"
    }

    cdl_interface CYGINT_HAL_ARM_AT91_SYS_INTERRUPT {
        display     "AT91 core has multiplexed system interrupts"    
        description "
            Some AT91 cores have a system controller which multiplexes
            many interrupts onto the system interrupt. When this interface
            is enabled the variant hal will perform a second level
            expansion of these interrupts"
    }

    cdl_interface CYGINT_HAL_ARM_AT91_PIT_HW {
        display     "Platform has a Periodic Interval Timer"
        description "
            This interface if implemented by HALs for CPU cores which
            have the Periodic Interval Timer."
    }

    cdl_option CYGBLD_HAL_ARM_AT91_TIMER_TC {
        display       "Use Timer Counter for eCos Clock"
        flavor        bool
        default_value 1
        requires      !CYGBLD_HAL_ARM_AT91_TIMER_PIT
        compile       timer_tc.c
        description   "
            Use a Timer Counter Channel to generate the eCos Clock."
    }

    cdl_option CYGBLD_HAL_ARM_AT91_TIMER_PIT {
        display       "Use Periodic Interval Timer for eCos Clock"
        flavor        bool
        default_value !CYGBLD_HAL_ARM_AT91_TIMER_TC
        requires      !CYGBLD_HAL_ARM_AT91_TIMER_TC
        active_if     CYGINT_HAL_ARM_AT91_PIT_HW
        compile       timer_pit.c
        description   "
            Use Periodic Interval Timer to generate the eCos Clock."
    }

    cdl_interface CYGINT_HAL_ARM_AT91_SERIAL_DBG_HW {
        display     "Platform has the DBG serial port"
        description "
            Some variants of the AT91 have a dedicated debug serial
            port. The HALs of such a variant should implement this interface
            so allowing the serial driver to the compiled"
    }

    cdl_option CYGBLD_HAL_ARM_AT91_SERIAL_DBG {
        display       "Enable the use of the DBG serial port"
        flavor        bool
        active_if     CYGINT_HAL_ARM_AT91_SERIAL_DBG_HW
        active_if     !CYGBLD_HAL_ARM_AT91_SERIAL_UART
        requires      CYGINT_HAL_ARM_AT91_SYS_INTERRUPT
        default_value 1

        compile       hal_diag_dbg.c 
        requires      CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL == 0
        requires      CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL == 0

        description   "
            The driver for the dedicated DBG UART will be compiled in the
            variant HAL when this option is enabled."
    }

    cdl_option CYGBLD_HAL_ARM_AT91_SERIAL_UART {
        display       "Enable the use of the UARTS for debug output"
        flavor        bool
        default_value 1
        compile       hal_diag.c 
        requires      !CYGBLD_HAL_ARM_AT91_SERIAL_DBG
        description   "        
            The driver for using the UARTS will be compiled in the
            variant HAL when this option is enabled."
    }

    cdl_component CYGBLD_HAL_ARM_AT91_DCC {
        display       "Enable the use of the DCC for debug output"
        flavor        bool
        default_value 0
        compile       hal_diag_dcc.c
        description   "
            A <serial> driver will be compiled and inserted into the
            vector table which does I/O via the DCC. The DCC is part of
            the JTAG interface and some JTAG devices made this interface
            available via telnet etc."
        
        cdl_option CYGBLD_HAL_ARM_AT91_DCC_CHANNEL {   
            display       "Channel the DCC port should use in the VV table"
            flavor        data
            default_value 2
            description   "
                The DCC driver has to be registered in the VV table of
                drivers. This option determines which entry in the
                table it will take. The default value will overwride
                the first serial port. "
        }
    }

    cdl_option CYGFUN_HAL_ARM_AT91_PROFILE_TIMER {
        display       "Use TC1 for gprof profiling"
        active_if     CYGPKG_PROFILE_GPROF
        flavor        bool
        default_value 1
        requires      !CYGPKG_HAL_ARM_AT91_JTST
        implements    CYGINT_PROFILE_HAL_TIMER
        description   "
            The AT91 variant HAL can provide support for gprof-based
            profiling. This uses timer TC1 to generate regular interrupts,
            and the interrupt handler records the PC at the time of the
            interrupt. However, TC1 is unavailable for this purpose on
            the JTST platform. Disable this option if you wish to provide
            an alternative profiling timer implementation."
    }
}
